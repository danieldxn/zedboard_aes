library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_package.BYTE;

entity multiply_2 is
	port (i : in BYTE;
			o : out BYTE
			);		
end multiply_2;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_package.BYTE;
entity multiply_3 is
	port (i : in BYTE;
			o : out BYTE
			);	
end multiply_3;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_package.BYTE;
entity multiply_9 is
	port (i : in BYTE;
			o : out BYTE
			);
end multiply_9;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_package.BYTE;
entity multiply_b is
	port (i : in BYTE;
			o : out BYTE
			);
end multiply_b;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_package.BYTE;
entity multiply_d is
	port (i : in BYTE;
			o : out BYTE
			);
end multiply_d;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_package.BYTE;
entity multiply_e is
	port (i : in std_logic_vector (7 downto 0); --This should be BYTE
			o : out std_logic_vector (7 downto 0) -- This should be BYTE
			);
end multiply_e;

architecture Behavioral of multiply_2 is

begin
	with i select o <=
		x"00" when x"00",
		x"02" when x"01",
		x"04" when x"02",
		x"06" when x"03",
		x"08" when x"04",
		x"0A" when x"05",
		x"0C" when x"06",
		x"0E" when x"07",
		x"10" when x"08",
		x"12" when x"09",
		x"14" when x"0A",
		x"16" when x"0B",
		x"18" when x"0C",
		x"1A" when x"0D",
		x"1C" when x"0E",
		x"1E" when x"0F",
		x"20" when x"10",
		x"22" when x"11",
		x"24" when x"12",
		x"26" when x"13",
		x"28" when x"14",
		x"2A" when x"15",
		x"2C" when x"16",
		x"2E" when x"17",
		x"30" when x"18",
		x"32" when x"19",
		x"34" when x"1A",
		x"36" when x"1B",
		x"38" when x"1C",
		x"3A" when x"1D",
		x"3C" when x"1E",
		x"3E" when x"1F",
		x"40" when x"20",
		x"42" when x"21",
		x"44" when x"22",
		x"46" when x"23",
		x"48" when x"24",
		x"4A" when x"25",
		x"4C" when x"26",
		x"4E" when x"27",
		x"50" when x"28",
		x"52" when x"29",
		x"54" when x"2A",
		x"56" when x"2B",
		x"58" when x"2C",
		x"5A" when x"2D",
		x"5C" when x"2E",
		x"5E" when x"2F",
		x"60" when x"30",
		x"62" when x"31",
		x"64" when x"32",
		x"66" when x"33",
		x"68" when x"34",
		x"6A" when x"35",
		x"6C" when x"36",
		x"6E" when x"37",
		x"70" when x"38",
		x"72" when x"39",
		x"74" when x"3A",
		x"76" when x"3B",
		x"78" when x"3C",
		x"7A" when x"3D",
		x"7C" when x"3E",
		x"7E" when x"3F",
		x"80" when x"40",
		x"82" when x"41",
		x"84" when x"42",
		x"86" when x"43",
		x"88" when x"44",
		x"8A" when x"45",
		x"8C" when x"46",
		x"8E" when x"47",
		x"90" when x"48",
		x"92" when x"49",
		x"94" when x"4A",
		x"96" when x"4B",
		x"98" when x"4C",
		x"9A" when x"4D",
		x"9C" when x"4E",
		x"9E" when x"4F",
		x"A0" when x"50",
		x"A2" when x"51",
		x"A4" when x"52",
		x"A6" when x"53",
		x"A8" when x"54",
		x"AA" when x"55",
		x"AC" when x"56",
		x"AE" when x"57",
		x"B0" when x"58",
		x"B2" when x"59",
		x"B4" when x"5A",
		x"B6" when x"5B",
		x"B8" when x"5C",
		x"BA" when x"5D",
		x"BC" when x"5E",
		x"BE" when x"5F",
		x"C0" when x"60",
		x"C2" when x"61",
		x"C4" when x"62",
		x"C6" when x"63",
		x"C8" when x"64",
		x"CA" when x"65",
		x"CC" when x"66",
		x"CE" when x"67",
		x"D0" when x"68",
		x"D2" when x"69",
		x"D4" when x"6A",
		x"D6" when x"6B",
		x"D8" when x"6C",
		x"DA" when x"6D",
		x"DC" when x"6E",
		x"DE" when x"6F",
		x"E0" when x"70",
		x"E2" when x"71",
		x"E4" when x"72",
		x"E6" when x"73",
		x"E8" when x"74",
		x"EA" when x"75",
		x"EC" when x"76",
		x"EE" when x"77",
		x"F0" when x"78",
		x"F2" when x"79",
		x"F4" when x"7A",
		x"F6" when x"7B",
		x"F8" when x"7C",
		x"FA" when x"7D",
		x"FC" when x"7E",
		x"FE" when x"7F",
		x"1B" when x"80",
		x"19" when x"81",
		x"1F" when x"82",
		x"1D" when x"83",
		x"13" when x"84",
		x"11" when x"85",
		x"17" when x"86",
		x"15" when x"87",
		x"0B" when x"88",
		x"09" when x"89",
		x"0F" when x"8A",
		x"0D" when x"8B",
		x"03" when x"8C",
		x"01" when x"8D",
		x"07" when x"8E",
		x"05" when x"8F",
		x"3B" when x"90",
		x"39" when x"91",
		x"3F" when x"92",
		x"3D" when x"93",
		x"33" when x"94",
		x"31" when x"95",
		x"37" when x"96",
		x"35" when x"97",
		x"2B" when x"98",
		x"29" when x"99",
		x"2F" when x"9A",
		x"2D" when x"9B",
		x"23" when x"9C",
		x"21" when x"9D",
		x"27" when x"9E",
		x"25" when x"9F",
		x"5B" when x"A0",
		x"59" when x"A1",
		x"5F" when x"A2",
		x"5D" when x"A3",
		x"53" when x"A4",
		x"51" when x"A5",
		x"57" when x"A6",
		x"55" when x"A7",
		x"4B" when x"A8",
		x"49" when x"A9",
		x"4F" when x"AA",
		x"4D" when x"AB",
		x"43" when x"AC",
		x"41" when x"AD",
		x"47" when x"AE",
		x"45" when x"AF",
		x"7B" when x"B0",
		x"79" when x"B1",
		x"7F" when x"B2",
		x"7D" when x"B3",
		x"73" when x"B4",
		x"71" when x"B5",
		x"77" when x"B6",
		x"75" when x"B7",
		x"6B" when x"B8",
		x"69" when x"B9",
		x"6F" when x"BA",
		x"6D" when x"BB",
		x"63" when x"BC",
		x"61" when x"BD",
		x"67" when x"BE",
		x"65" when x"BF",
		x"9B" when x"C0",
		x"99" when x"C1",
		x"9F" when x"C2",
		x"9D" when x"C3",
		x"93" when x"C4",
		x"91" when x"C5",
		x"97" when x"C6",
		x"95" when x"C7",
		x"8B" when x"C8",
		x"89" when x"C9",
		x"8F" when x"CA",
		x"8D" when x"CB",
		x"83" when x"CC",
		x"81" when x"CD",
		x"87" when x"CE",
		x"85" when x"CF",
		x"BB" when x"D0",
		x"B9" when x"D1",
		x"BF" when x"D2",
		x"BD" when x"D3",
		x"B3" when x"D4",
		x"B1" when x"D5",
		x"B7" when x"D6",
		x"B5" when x"D7",
		x"AB" when x"D8",
		x"A9" when x"D9",
		x"AF" when x"DA",
		x"AD" when x"DB",
		x"A3" when x"DC",
		x"A1" when x"DD",
		x"A7" when x"DE",
		x"A5" when x"DF",
		x"DB" when x"E0",
		x"D9" when x"E1",
		x"DF" when x"E2",
		x"DD" when x"E3",
		x"D3" when x"E4",
		x"D1" when x"E5",
		x"D7" when x"E6",
		x"D5" when x"E7",
		x"CB" when x"E8",
		x"C9" when x"E9",
		x"CF" when x"EA",
		x"CD" when x"EB",
		x"C3" when x"EC",
		x"C1" when x"ED",
		x"C7" when x"EE",
		x"C5" when x"EF",
		x"FB" when x"F0",
		x"F9" when x"F1",
		x"FF" when x"F2",
		x"FD" when x"F3",
		x"F3" when x"F4",
		x"F1" when x"F5",
		x"F7" when x"F6",
		x"F5" when x"F7",
		x"EB" when x"F8",
		x"E9" when x"F9",
		x"EF" when x"FA",
		x"ED" when x"FB",
		x"E3" when x"FC",
		x"E1" when x"FD",
		x"E7" when x"FE",
		x"E5" when x"FF",
		x"00" when others;

end Behavioral;

architecture Behavioral of multiply_3 is

begin
	with i select o <=
		x"00" when x"00",
		x"03" when x"01",
		x"06" when x"02",
		x"05" when x"03",
		x"0C" when x"04",
		x"0F" when x"05",
		x"0A" when x"06",
		x"09" when x"07",
		x"18" when x"08",
		x"1B" when x"09",
		x"1E" when x"0A",
		x"1D" when x"0B",
		x"14" when x"0C",
		x"17" when x"0D",
		x"12" when x"0E",
		x"11" when x"0F",
		x"30" when x"10",
		x"33" when x"11",
		x"36" when x"12",
		x"35" when x"13",
		x"3C" when x"14",
		x"3F" when x"15",
		x"3A" when x"16",
		x"39" when x"17",
		x"28" when x"18",
		x"2B" when x"19",
		x"2E" when x"1A",
		x"2D" when x"1B",
		x"24" when x"1C",
		x"27" when x"1D",
		x"22" when x"1E",
		x"21" when x"1F",
		x"60" when x"20",
		x"63" when x"21",
		x"66" when x"22",
		x"65" when x"23",
		x"6C" when x"24",
		x"6F" when x"25",
		x"6A" when x"26",
		x"69" when x"27",
		x"78" when x"28",
		x"7B" when x"29",
		x"7E" when x"2A",
		x"7D" when x"2B",
		x"74" when x"2C",
		x"77" when x"2D",
		x"72" when x"2E",
		x"71" when x"2F",
		x"50" when x"30",
		x"53" when x"31",
		x"56" when x"32",
		x"55" when x"33",
		x"5C" when x"34",
		x"5F" when x"35",
		x"5A" when x"36",
		x"59" when x"37",
		x"48" when x"38",
		x"4B" when x"39",
		x"4E" when x"3A",
		x"4D" when x"3B",
		x"44" when x"3C",
		x"47" when x"3D",
		x"42" when x"3E",
		x"41" when x"3F",
		x"C0" when x"40",
		x"C3" when x"41",
		x"C6" when x"42",
		x"C5" when x"43",
		x"CC" when x"44",
		x"CF" when x"45",
		x"CA" when x"46",
		x"C9" when x"47",
		x"D8" when x"48",
		x"DB" when x"49",
		x"DE" when x"4A",
		x"DD" when x"4B",
		x"D4" when x"4C",
		x"D7" when x"4D",
		x"D2" when x"4E",
		x"D1" when x"4F",
		x"F0" when x"50",
		x"F3" when x"51",
		x"F6" when x"52",
		x"F5" when x"53",
		x"FC" when x"54",
		x"FF" when x"55",
		x"FA" when x"56",
		x"F9" when x"57",
		x"E8" when x"58",
		x"EB" when x"59",
		x"EE" when x"5A",
		x"ED" when x"5B",
		x"E4" when x"5C",
		x"E7" when x"5D",
		x"E2" when x"5E",
		x"E1" when x"5F",
		x"A0" when x"60",
		x"A3" when x"61",
		x"A6" when x"62",
		x"A5" when x"63",
		x"AC" when x"64",
		x"AF" when x"65",
		x"AA" when x"66",
		x"A9" when x"67",
		x"B8" when x"68",
		x"BB" when x"69",
		x"BE" when x"6A",
		x"BD" when x"6B",
		x"B4" when x"6C",
		x"B7" when x"6D",
		x"B2" when x"6E",
		x"B1" when x"6F",
		x"90" when x"70",
		x"93" when x"71",
		x"96" when x"72",
		x"95" when x"73",
		x"9C" when x"74",
		x"9F" when x"75",
		x"9A" when x"76",
		x"99" when x"77",
		x"88" when x"78",
		x"8B" when x"79",
		x"8E" when x"7A",
		x"8D" when x"7B",
		x"84" when x"7C",
		x"87" when x"7D",
		x"82" when x"7E",
		x"81" when x"7F",
		x"9B" when x"80",
		x"98" when x"81",
		x"9D" when x"82",
		x"9E" when x"83",
		x"97" when x"84",
		x"94" when x"85",
		x"91" when x"86",
		x"92" when x"87",
		x"83" when x"88",
		x"80" when x"89",
		x"85" when x"8A",
		x"86" when x"8B",
		x"8F" when x"8C",
		x"8C" when x"8D",
		x"89" when x"8E",
		x"8A" when x"8F",
		x"AB" when x"90",
		x"A8" when x"91",
		x"AD" when x"92",
		x"AE" when x"93",
		x"A7" when x"94",
		x"A4" when x"95",
		x"A1" when x"96",
		x"A2" when x"97",
		x"B3" when x"98",
		x"B0" when x"99",
		x"B5" when x"9A",
		x"B6" when x"9B",
		x"BF" when x"9C",
		x"BC" when x"9D",
		x"B9" when x"9E",
		x"BA" when x"9F",
		x"FB" when x"A0",
		x"F8" when x"A1",
		x"FD" when x"A2",
		x"FE" when x"A3",
		x"F7" when x"A4",
		x"F4" when x"A5",
		x"F1" when x"A6",
		x"F2" when x"A7",
		x"E3" when x"A8",
		x"E0" when x"A9",
		x"E5" when x"AA",
		x"E6" when x"AB",
		x"EF" when x"AC",
		x"EC" when x"AD",
		x"E9" when x"AE",
		x"EA" when x"AF",
		x"CB" when x"B0",
		x"C8" when x"B1",
		x"CD" when x"B2",
		x"CE" when x"B3",
		x"C7" when x"B4",
		x"C4" when x"B5",
		x"C1" when x"B6",
		x"C2" when x"B7",
		x"D3" when x"B8",
		x"D0" when x"B9",
		x"D5" when x"BA",
		x"D6" when x"BB",
		x"DF" when x"BC",
		x"DC" when x"BD",
		x"D9" when x"BE",
		x"DA" when x"BF",
		x"5B" when x"C0",
		x"58" when x"C1",
		x"5D" when x"C2",
		x"5E" when x"C3",
		x"57" when x"C4",
		x"54" when x"C5",
		x"51" when x"C6",
		x"52" when x"C7",
		x"43" when x"C8",
		x"40" when x"C9",
		x"45" when x"CA",
		x"46" when x"CB",
		x"4F" when x"CC",
		x"4C" when x"CD",
		x"49" when x"CE",
		x"4A" when x"CF",
		x"6B" when x"D0",
		x"68" when x"D1",
		x"6D" when x"D2",
		x"6E" when x"D3",
		x"67" when x"D4",
		x"64" when x"D5",
		x"61" when x"D6",
		x"62" when x"D7",
		x"73" when x"D8",
		x"70" when x"D9",
		x"75" when x"DA",
		x"76" when x"DB",
		x"7F" when x"DC",
		x"7C" when x"DD",
		x"79" when x"DE",
		x"7A" when x"DF",
		x"3B" when x"E0",
		x"38" when x"E1",
		x"3D" when x"E2",
		x"3E" when x"E3",
		x"37" when x"E4",
		x"34" when x"E5",
		x"31" when x"E6",
		x"32" when x"E7",
		x"23" when x"E8",
		x"20" when x"E9",
		x"25" when x"EA",
		x"26" when x"EB",
		x"2F" when x"EC",
		x"2C" when x"ED",
		x"29" when x"EE",
		x"2A" when x"EF",
		x"0B" when x"F0",
		x"08" when x"F1",
		x"0D" when x"F2",
		x"0E" when x"F3",
		x"07" when x"F4",
		x"04" when x"F5",
		x"01" when x"F6",
		x"02" when x"F7",
		x"13" when x"F8",
		x"10" when x"F9",
		x"15" when x"FA",
		x"16" when x"FB",
		x"1F" when x"FC",
		x"1C" when x"FD",
		x"19" when x"FE",
		x"1A" when x"FF",
		x"00" when others;

end Behavioral;

architecture Behavioral of multiply_9 is

begin
	with i select o <=
		x"00" when x"00",
		x"09" when x"01",
		x"12" when x"02",
		x"1B" when x"03",
		x"24" when x"04",
		x"2D" when x"05",
		x"36" when x"06",
		x"3F" when x"07",
		x"48" when x"08",
		x"41" when x"09",
		x"5A" when x"0A",
		x"53" when x"0B",
		x"6C" when x"0C",
		x"65" when x"0D",
		x"7E" when x"0E",
		x"77" when x"0F",
		x"90" when x"10",
		x"99" when x"11",
		x"82" when x"12",
		x"8B" when x"13",
		x"B4" when x"14",
		x"BD" when x"15",
		x"A6" when x"16",
		x"AF" when x"17",
		x"D8" when x"18",
		x"D1" when x"19",
		x"CA" when x"1A",
		x"C3" when x"1B",
		x"FC" when x"1C",
		x"F5" when x"1D",
		x"EE" when x"1E",
		x"E7" when x"1F",
		x"3B" when x"20",
		x"32" when x"21",
		x"29" when x"22",
		x"20" when x"23",
		x"1F" when x"24",
		x"16" when x"25",
		x"0D" when x"26",
		x"04" when x"27",
		x"73" when x"28",
		x"7A" when x"29",
		x"61" when x"2A",
		x"68" when x"2B",
		x"57" when x"2C",
		x"5E" when x"2D",
		x"45" when x"2E",
		x"4C" when x"2F",
		x"AB" when x"30",
		x"A2" when x"31",
		x"B9" when x"32",
		x"B0" when x"33",
		x"8F" when x"34",
		x"86" when x"35",
		x"9D" when x"36",
		x"94" when x"37",
		x"E3" when x"38",
		x"EA" when x"39",
		x"F1" when x"3A",
		x"F8" when x"3B",
		x"C7" when x"3C",
		x"CE" when x"3D",
		x"D5" when x"3E",
		x"DC" when x"3F",
		x"76" when x"40",
		x"7F" when x"41",
		x"64" when x"42",
		x"6D" when x"43",
		x"52" when x"44",
		x"5B" when x"45",
		x"40" when x"46",
		x"49" when x"47",
		x"3E" when x"48",
		x"37" when x"49",
		x"2C" when x"4A",
		x"25" when x"4B",
		x"1A" when x"4C",
		x"13" when x"4D",
		x"08" when x"4E",
		x"01" when x"4F",
		x"E6" when x"50",
		x"EF" when x"51",
		x"F4" when x"52",
		x"FD" when x"53",
		x"C2" when x"54",
		x"CB" when x"55",
		x"D0" when x"56",
		x"D9" when x"57",
		x"AE" when x"58",
		x"A7" when x"59",
		x"BC" when x"5A",
		x"B5" when x"5B",
		x"8A" when x"5C",
		x"83" when x"5D",
		x"98" when x"5E",
		x"91" when x"5F",
		x"4D" when x"60",
		x"44" when x"61",
		x"5F" when x"62",
		x"56" when x"63",
		x"69" when x"64",
		x"60" when x"65",
		x"7B" when x"66",
		x"72" when x"67",
		x"05" when x"68",
		x"0C" when x"69",
		x"17" when x"6A",
		x"1E" when x"6B",
		x"21" when x"6C",
		x"28" when x"6D",
		x"33" when x"6E",
		x"3A" when x"6F",
		x"DD" when x"70",
		x"D4" when x"71",
		x"CF" when x"72",
		x"C6" when x"73",
		x"F9" when x"74",
		x"F0" when x"75",
		x"EB" when x"76",
		x"E2" when x"77",
		x"95" when x"78",
		x"9C" when x"79",
		x"87" when x"7A",
		x"8E" when x"7B",
		x"B1" when x"7C",
		x"B8" when x"7D",
		x"A3" when x"7E",
		x"AA" when x"7F",
		x"EC" when x"80",
		x"E5" when x"81",
		x"FE" when x"82",
		x"F7" when x"83",
		x"C8" when x"84",
		x"C1" when x"85",
		x"DA" when x"86",
		x"D3" when x"87",
		x"A4" when x"88",
		x"AD" when x"89",
		x"B6" when x"8A",
		x"BF" when x"8B",
		x"80" when x"8C",
		x"89" when x"8D",
		x"92" when x"8E",
		x"9B" when x"8F",
		x"7C" when x"90",
		x"75" when x"91",
		x"6E" when x"92",
		x"67" when x"93",
		x"58" when x"94",
		x"51" when x"95",
		x"4A" when x"96",
		x"43" when x"97",
		x"34" when x"98",
		x"3D" when x"99",
		x"26" when x"9A",
		x"2F" when x"9B",
		x"10" when x"9C",
		x"19" when x"9D",
		x"02" when x"9E",
		x"0B" when x"9F",
		x"D7" when x"A0",
		x"DE" when x"A1",
		x"C5" when x"A2",
		x"CC" when x"A3",
		x"F3" when x"A4",
		x"FA" when x"A5",
		x"E1" when x"A6",
		x"E8" when x"A7",
		x"9F" when x"A8",
		x"96" when x"A9",
		x"8D" when x"AA",
		x"84" when x"AB",
		x"BB" when x"AC",
		x"B2" when x"AD",
		x"A9" when x"AE",
		x"A0" when x"AF",
		x"47" when x"B0",
		x"4E" when x"B1",
		x"55" when x"B2",
		x"5C" when x"B3",
		x"63" when x"B4",
		x"6A" when x"B5",
		x"71" when x"B6",
		x"78" when x"B7",
		x"0F" when x"B8",
		x"06" when x"B9",
		x"1D" when x"BA",
		x"14" when x"BB",
		x"2B" when x"BC",
		x"22" when x"BD",
		x"39" when x"BE",
		x"30" when x"BF",
		x"9A" when x"C0",
		x"93" when x"C1",
		x"88" when x"C2",
		x"81" when x"C3",
		x"BE" when x"C4",
		x"B7" when x"C5",
		x"AC" when x"C6",
		x"A5" when x"C7",
		x"D2" when x"C8",
		x"DB" when x"C9",
		x"C0" when x"CA",
		x"C9" when x"CB",
		x"F6" when x"CC",
		x"FF" when x"CD",
		x"E4" when x"CE",
		x"ED" when x"CF",
		x"0A" when x"D0",
		x"03" when x"D1",
		x"18" when x"D2",
		x"11" when x"D3",
		x"2E" when x"D4",
		x"27" when x"D5",
		x"3C" when x"D6",
		x"35" when x"D7",
		x"42" when x"D8",
		x"4B" when x"D9",
		x"50" when x"DA",
		x"59" when x"DB",
		x"66" when x"DC",
		x"6F" when x"DD",
		x"74" when x"DE",
		x"7D" when x"DF",
		x"A1" when x"E0",
		x"A8" when x"E1",
		x"B3" when x"E2",
		x"BA" when x"E3",
		x"85" when x"E4",
		x"8C" when x"E5",
		x"97" when x"E6",
		x"9E" when x"E7",
		x"E9" when x"E8",
		x"E0" when x"E9",
		x"FB" when x"EA",
		x"F2" when x"EB",
		x"CD" when x"EC",
		x"C4" when x"ED",
		x"DF" when x"EE",
		x"D6" when x"EF",
		x"31" when x"F0",
		x"38" when x"F1",
		x"23" when x"F2",
		x"2A" when x"F3",
		x"15" when x"F4",
		x"1C" when x"F5",
		x"07" when x"F6",
		x"0E" when x"F7",
		x"79" when x"F8",
		x"70" when x"F9",
		x"6B" when x"FA",
		x"62" when x"FB",
		x"5D" when x"FC",
		x"54" when x"FD",
		x"4F" when x"FE",
		x"46" when x"FF",
		x"00" when others;  

end Behavioral;

architecture Behavioral of multiply_b is

begin
	with i select o <=
		x"00" when x"00",
		x"0B" when x"01",
		x"16" when x"02",
		x"1D" when x"03",
		x"2C" when x"04",
		x"27" when x"05",
		x"3A" when x"06",
		x"31" when x"07",
		x"58" when x"08",
		x"53" when x"09",
		x"4E" when x"0A",
		x"45" when x"0B",
		x"74" when x"0C",
		x"7F" when x"0D",
		x"62" when x"0E",
		x"69" when x"0F",
		x"B0" when x"10",
		x"BB" when x"11",
		x"A6" when x"12",
		x"AD" when x"13",
		x"9C" when x"14",
		x"97" when x"15",
		x"8A" when x"16",
		x"81" when x"17",
		x"E8" when x"18",
		x"E3" when x"19",
		x"FE" when x"1A",
		x"F5" when x"1B",
		x"C4" when x"1C",
		x"CF" when x"1D",
		x"D2" when x"1E",
		x"D9" when x"1F",
		x"7B" when x"20",
		x"70" when x"21",
		x"6D" when x"22",
		x"66" when x"23",
		x"57" when x"24",
		x"5C" when x"25",
		x"41" when x"26",
		x"4A" when x"27",
		x"23" when x"28",
		x"28" when x"29",
		x"35" when x"2A",
		x"3E" when x"2B",
		x"0F" when x"2C",
		x"04" when x"2D",
		x"19" when x"2E",
		x"12" when x"2F",
		x"CB" when x"30",
		x"C0" when x"31",
		x"DD" when x"32",
		x"D6" when x"33",
		x"E7" when x"34",
		x"EC" when x"35",
		x"F1" when x"36",
		x"FA" when x"37",
		x"93" when x"38",
		x"98" when x"39",
		x"85" when x"3A",
		x"8E" when x"3B",
		x"BF" when x"3C",
		x"B4" when x"3D",
		x"A9" when x"3E",
		x"A2" when x"3F",
		x"F6" when x"40",
		x"FD" when x"41",
		x"E0" when x"42",
		x"EB" when x"43",
		x"DA" when x"44",
		x"D1" when x"45",
		x"CC" when x"46",
		x"C7" when x"47",
		x"AE" when x"48",
		x"A5" when x"49",
		x"B8" when x"4A",
		x"B3" when x"4B",
		x"82" when x"4C",
		x"89" when x"4D",
		x"94" when x"4E",
		x"9F" when x"4F",
		x"46" when x"50",
		x"4D" when x"51",
		x"50" when x"52",
		x"5B" when x"53",
		x"6A" when x"54",
		x"61" when x"55",
		x"7C" when x"56",
		x"77" when x"57",
		x"1E" when x"58",
		x"15" when x"59",
		x"08" when x"5A",
		x"03" when x"5B",
		x"32" when x"5C",
		x"39" when x"5D",
		x"24" when x"5E",
		x"2F" when x"5F",
		x"8D" when x"60",
		x"86" when x"61",
		x"9B" when x"62",
		x"90" when x"63",
		x"A1" when x"64",
		x"AA" when x"65",
		x"B7" when x"66",
		x"BC" when x"67",
		x"D5" when x"68",
		x"DE" when x"69",
		x"C3" when x"6A",
		x"C8" when x"6B",
		x"F9" when x"6C",
		x"F2" when x"6D",
		x"EF" when x"6E",
		x"E4" when x"6F",
		x"3D" when x"70",
		x"36" when x"71",
		x"2B" when x"72",
		x"20" when x"73",
		x"11" when x"74",
		x"1A" when x"75",
		x"07" when x"76",
		x"0C" when x"77",
		x"65" when x"78",
		x"6E" when x"79",
		x"73" when x"7A",
		x"78" when x"7B",
		x"49" when x"7C",
		x"42" when x"7D",
		x"5F" when x"7E",
		x"54" when x"7F",
		x"F7" when x"80",
		x"FC" when x"81",
		x"E1" when x"82",
		x"EA" when x"83",
		x"DB" when x"84",
		x"D0" when x"85",
		x"CD" when x"86",
		x"C6" when x"87",
		x"AF" when x"88",
		x"A4" when x"89",
		x"B9" when x"8A",
		x"B2" when x"8B",
		x"83" when x"8C",
		x"88" when x"8D",
		x"95" when x"8E",
		x"9E" when x"8F",
		x"47" when x"90",
		x"4C" when x"91",
		x"51" when x"92",
		x"5A" when x"93",
		x"6B" when x"94",
		x"60" when x"95",
		x"7D" when x"96",
		x"76" when x"97",
		x"1F" when x"98",
		x"14" when x"99",
		x"09" when x"9A",
		x"02" when x"9B",
		x"33" when x"9C",
		x"38" when x"9D",
		x"25" when x"9E",
		x"2E" when x"9F",
		x"8C" when x"A0",
		x"87" when x"A1",
		x"9A" when x"A2",
		x"91" when x"A3",
		x"A0" when x"A4",
		x"AB" when x"A5",
		x"B6" when x"A6",
		x"BD" when x"A7",
		x"D4" when x"A8",
		x"DF" when x"A9",
		x"C2" when x"AA",
		x"C9" when x"AB",
		x"F8" when x"AC",
		x"F3" when x"AD",
		x"EE" when x"AE",
		x"E5" when x"AF",
		x"3C" when x"B0",
		x"37" when x"B1",
		x"2A" when x"B2",
		x"21" when x"B3",
		x"10" when x"B4",
		x"1B" when x"B5",
		x"06" when x"B6",
		x"0D" when x"B7",
		x"64" when x"B8",
		x"6F" when x"B9",
		x"72" when x"BA",
		x"79" when x"BB",
		x"48" when x"BC",
		x"43" when x"BD",
		x"5E" when x"BE",
		x"55" when x"BF",
		x"01" when x"C0",
		x"0A" when x"C1",
		x"17" when x"C2",
		x"1C" when x"C3",
		x"2D" when x"C4",
		x"26" when x"C5",
		x"3B" when x"C6",
		x"30" when x"C7",
		x"59" when x"C8",
		x"52" when x"C9",
		x"4F" when x"CA",
		x"44" when x"CB",
		x"75" when x"CC",
		x"7E" when x"CD",
		x"63" when x"CE",
		x"68" when x"CF",
		x"B1" when x"D0",
		x"BA" when x"D1",
		x"A7" when x"D2",
		x"AC" when x"D3",
		x"9D" when x"D4",
		x"96" when x"D5",
		x"8B" when x"D6",
		x"80" when x"D7",
		x"E9" when x"D8",
		x"E2" when x"D9",
		x"FF" when x"DA",
		x"F4" when x"DB",
		x"C5" when x"DC",
		x"CE" when x"DD",
		x"D3" when x"DE",
		x"D8" when x"DF",
		x"7A" when x"E0",
		x"71" when x"E1",
		x"6C" when x"E2",
		x"67" when x"E3",
		x"56" when x"E4",
		x"5D" when x"E5",
		x"40" when x"E6",
		x"4B" when x"E7",
		x"22" when x"E8",
		x"29" when x"E9",
		x"34" when x"EA",
		x"3F" when x"EB",
		x"0E" when x"EC",
		x"05" when x"ED",
		x"18" when x"EE",
		x"13" when x"EF",
		x"CA" when x"F0",
		x"C1" when x"F1",
		x"DC" when x"F2",
		x"D7" when x"F3",
		x"E6" when x"F4",
		x"ED" when x"F5",
		x"F0" when x"F6",
		x"FB" when x"F7",
		x"92" when x"F8",
		x"99" when x"F9",
		x"84" when x"FA",
		x"8F" when x"FB",
		x"BE" when x"FC",
		x"B5" when x"FD",
		x"A8" when x"FE",
		x"A3" when x"FF",
		x"00" when others;

end Behavioral;

architecture Behavioral of multiply_d is

begin
	with i select o <=
		x"00" when x"00",
		x"0D" when x"01",
		x"1A" when x"02",
		x"17" when x"03",
		x"34" when x"04",
		x"39" when x"05",
		x"2E" when x"06",
		x"23" when x"07",
		x"68" when x"08",
		x"65" when x"09",
		x"72" when x"0A",
		x"7F" when x"0B",
		x"5C" when x"0C",
		x"51" when x"0D",
		x"46" when x"0E",
		x"4B" when x"0F",
		x"D0" when x"10",
		x"DD" when x"11",
		x"CA" when x"12",
		x"C7" when x"13",
		x"E4" when x"14",
		x"E9" when x"15",
		x"FE" when x"16",
		x"F3" when x"17",
		x"B8" when x"18",
		x"B5" when x"19",
		x"A2" when x"1A",
		x"AF" when x"1B",
		x"8C" when x"1C",
		x"81" when x"1D",
		x"96" when x"1E",
		x"9B" when x"1F",
		x"BB" when x"20",
		x"B6" when x"21",
		x"A1" when x"22",
		x"AC" when x"23",
		x"8F" when x"24",
		x"82" when x"25",
		x"95" when x"26",
		x"98" when x"27",
		x"D3" when x"28",
		x"DE" when x"29",
		x"C9" when x"2A",
		x"C4" when x"2B",
		x"E7" when x"2C",
		x"EA" when x"2D",
		x"FD" when x"2E",
		x"F0" when x"2F",
		x"6B" when x"30",
		x"66" when x"31",
		x"71" when x"32",
		x"7C" when x"33",
		x"5F" when x"34",
		x"52" when x"35",
		x"45" when x"36",
		x"48" when x"37",
		x"03" when x"38",
		x"0E" when x"39",
		x"19" when x"3A",
		x"14" when x"3B",
		x"37" when x"3C",
		x"3A" when x"3D",
		x"2D" when x"3E",
		x"20" when x"3F",
		x"6D" when x"40",
		x"60" when x"41",
		x"77" when x"42",
		x"7A" when x"43",
		x"59" when x"44",
		x"54" when x"45",
		x"43" when x"46",
		x"4E" when x"47",
		x"05" when x"48",
		x"08" when x"49",
		x"1F" when x"4A",
		x"12" when x"4B",
		x"31" when x"4C",
		x"3C" when x"4D",
		x"2B" when x"4E",
		x"26" when x"4F",
		x"BD" when x"50",
		x"B0" when x"51",
		x"A7" when x"52",
		x"AA" when x"53",
		x"89" when x"54",
		x"84" when x"55",
		x"93" when x"56",
		x"9E" when x"57",
		x"D5" when x"58",
		x"D8" when x"59",
		x"CF" when x"5A",
		x"C2" when x"5B",
		x"E1" when x"5C",
		x"EC" when x"5D",
		x"FB" when x"5E",
		x"F6" when x"5F",
		x"D6" when x"60",
		x"DB" when x"61",
		x"CC" when x"62",
		x"C1" when x"63",
		x"E2" when x"64",
		x"EF" when x"65",
		x"F8" when x"66",
		x"F5" when x"67",
		x"BE" when x"68",
		x"B3" when x"69",
		x"A4" when x"6A",
		x"A9" when x"6B",
		x"8A" when x"6C",
		x"87" when x"6D",
		x"90" when x"6E",
		x"9D" when x"6F",
		x"06" when x"70",
		x"0B" when x"71",
		x"1C" when x"72",
		x"11" when x"73",
		x"32" when x"74",
		x"3F" when x"75",
		x"28" when x"76",
		x"25" when x"77",
		x"6E" when x"78",
		x"63" when x"79",
		x"74" when x"7A",
		x"79" when x"7B",
		x"5A" when x"7C",
		x"57" when x"7D",
		x"40" when x"7E",
		x"4D" when x"7F",
		x"DA" when x"80",
		x"D7" when x"81",
		x"C0" when x"82",
		x"CD" when x"83",
		x"EE" when x"84",
		x"E3" when x"85",
		x"F4" when x"86",
		x"F9" when x"87",
		x"B2" when x"88",
		x"BF" when x"89",
		x"A8" when x"8A",
		x"A5" when x"8B",
		x"86" when x"8C",
		x"8B" when x"8D",
		x"9C" when x"8E",
		x"91" when x"8F",
		x"0A" when x"90",
		x"07" when x"91",
		x"10" when x"92",
		x"1D" when x"93",
		x"3E" when x"94",
		x"33" when x"95",
		x"24" when x"96",
		x"29" when x"97",
		x"62" when x"98",
		x"6F" when x"99",
		x"78" when x"9A",
		x"75" when x"9B",
		x"56" when x"9C",
		x"5B" when x"9D",
		x"4C" when x"9E",
		x"41" when x"9F",
		x"61" when x"A0",
		x"6C" when x"A1",
		x"7B" when x"A2",
		x"76" when x"A3",
		x"55" when x"A4",
		x"58" when x"A5",
		x"4F" when x"A6",
		x"42" when x"A7",
		x"09" when x"A8",
		x"04" when x"A9",
		x"13" when x"AA",
		x"1E" when x"AB",
		x"3D" when x"AC",
		x"30" when x"AD",
		x"27" when x"AE",
		x"2A" when x"AF",
		x"B1" when x"B0",
		x"BC" when x"B1",
		x"AB" when x"B2",
		x"A6" when x"B3",
		x"85" when x"B4",
		x"88" when x"B5",
		x"9F" when x"B6",
		x"92" when x"B7",
		x"D9" when x"B8",
		x"D4" when x"B9",
		x"C3" when x"BA",
		x"CE" when x"BB",
		x"ED" when x"BC",
		x"E0" when x"BD",
		x"F7" when x"BE",
		x"FA" when x"BF",
		x"B7" when x"C0",
		x"BA" when x"C1",
		x"AD" when x"C2",
		x"A0" when x"C3",
		x"83" when x"C4",
		x"8E" when x"C5",
		x"99" when x"C6",
		x"94" when x"C7",
		x"DF" when x"C8",
		x"D2" when x"C9",
		x"C5" when x"CA",
		x"C8" when x"CB",
		x"EB" when x"CC",
		x"E6" when x"CD",
		x"F1" when x"CE",
		x"FC" when x"CF",
		x"67" when x"D0",
		x"6A" when x"D1",
		x"7D" when x"D2",
		x"70" when x"D3",
		x"53" when x"D4",
		x"5E" when x"D5",
		x"49" when x"D6",
		x"44" when x"D7",
		x"0F" when x"D8",
		x"02" when x"D9",
		x"15" when x"DA",
		x"18" when x"DB",
		x"3B" when x"DC",
		x"36" when x"DD",
		x"21" when x"DE",
		x"2C" when x"DF",
		x"0C" when x"E0",
		x"01" when x"E1",
		x"16" when x"E2",
		x"1B" when x"E3",
		x"38" when x"E4",
		x"35" when x"E5",
		x"22" when x"E6",
		x"2F" when x"E7",
		x"64" when x"E8",
		x"69" when x"E9",
		x"7E" when x"EA",
		x"73" when x"EB",
		x"50" when x"EC",
		x"5D" when x"ED",
		x"4A" when x"EE",
		x"47" when x"EF",
		x"DC" when x"F0",
		x"D1" when x"F1",
		x"C6" when x"F2",
		x"CB" when x"F3",
		x"E8" when x"F4",
		x"E5" when x"F5",
		x"F2" when x"F6",
		x"FF" when x"F7",
		x"B4" when x"F8",
		x"B9" when x"F9",
		x"AE" when x"FA",
		x"A3" when x"FB",
		x"80" when x"FC",
		x"8D" when x"FD",
		x"9A" when x"FE",
		x"97" when x"FF",
		x"00" when others;

end Behavioral;

architecture Behavioral of multiply_e is
	
begin
	with i select o <=
		x"00" when x"00",
		x"0E" when x"01",
		x"1C" when x"02",
		x"12" when x"03",
		x"38" when x"04",
		x"36" when x"05",
		x"24" when x"06",
		x"2A" when x"07",
		x"70" when x"08",
		x"7E" when x"09",
		x"6C" when x"0A",
		x"62" when x"0B",
		x"48" when x"0C",
		x"46" when x"0D",
		x"54" when x"0E",
		x"5A" when x"0F",
		x"E0" when x"10",
		x"EE" when x"11",
		x"FC" when x"12",
		x"F2" when x"13",
		x"D8" when x"14",
		x"D6" when x"15",
		x"C4" when x"16",
		x"CA" when x"17",
		x"90" when x"18",
		x"9E" when x"19",
		x"8C" when x"1A",
		x"82" when x"1B",
		x"A8" when x"1C",
		x"A6" when x"1D",
		x"B4" when x"1E",
		x"BA" when x"1F",
		x"DB" when x"20",
		x"D5" when x"21",
		x"C7" when x"22",
		x"C9" when x"23",
		x"E3" when x"24",
		x"ED" when x"25",
		x"FF" when x"26",
		x"F1" when x"27",
		x"AB" when x"28",
		x"A5" when x"29",
		x"B7" when x"2A",
		x"B9" when x"2B",
		x"93" when x"2C",
		x"9D" when x"2D",
		x"8F" when x"2E",
		x"81" when x"2F",
		x"3B" when x"30",
		x"35" when x"31",
		x"27" when x"32",
		x"29" when x"33",
		x"03" when x"34",
		x"0D" when x"35",
		x"1F" when x"36",
		x"11" when x"37",
		x"4B" when x"38",
		x"45" when x"39",
		x"57" when x"3A",
		x"59" when x"3B",
		x"73" when x"3C",
		x"7D" when x"3D",
		x"6F" when x"3E",
		x"61" when x"3F",
		x"AD" when x"40",
		x"A3" when x"41",
		x"B1" when x"42",
		x"BF" when x"43",
		x"95" when x"44",
		x"9B" when x"45",
		x"89" when x"46",
		x"87" when x"47",
		x"DD" when x"48",
		x"D3" when x"49",
		x"C1" when x"4A",
		x"CF" when x"4B",
		x"E5" when x"4C",
		x"EB" when x"4D",
		x"F9" when x"4E",
		x"F7" when x"4F",
		x"4D" when x"50",
		x"43" when x"51",
		x"51" when x"52",
		x"5F" when x"53",
		x"75" when x"54",
		x"7B" when x"55",
		x"69" when x"56",
		x"67" when x"57",
		x"3D" when x"58",
		x"33" when x"59",
		x"21" when x"5A",
		x"2F" when x"5B",
		x"05" when x"5C",
		x"0B" when x"5D",
		x"19" when x"5E",
		x"17" when x"5F",
		x"76" when x"60",
		x"78" when x"61",
		x"6A" when x"62",
		x"64" when x"63",
		x"4E" when x"64",
		x"40" when x"65",
		x"52" when x"66",
		x"5C" when x"67",
		x"06" when x"68",
		x"08" when x"69",
		x"1A" when x"6A",
		x"14" when x"6B",
		x"3E" when x"6C",
		x"30" when x"6D",
		x"22" when x"6E",
		x"2C" when x"6F",
		x"96" when x"70",
		x"98" when x"71",
		x"8A" when x"72",
		x"84" when x"73",
		x"AE" when x"74",
		x"A0" when x"75",
		x"B2" when x"76",
		x"BC" when x"77",
		x"E6" when x"78",
		x"E8" when x"79",
		x"FA" when x"7A",
		x"F4" when x"7B",
		x"DE" when x"7C",
		x"D0" when x"7D",
		x"C2" when x"7E",
		x"CC" when x"7F",
		x"41" when x"80",
		x"4F" when x"81",
		x"5D" when x"82",
		x"53" when x"83",
		x"79" when x"84",
		x"77" when x"85",
		x"65" when x"86",
		x"6B" when x"87",
		x"31" when x"88",
		x"3F" when x"89",
		x"2D" when x"8A",
		x"23" when x"8B",
		x"09" when x"8C",
		x"07" when x"8D",
		x"15" when x"8E",
		x"1B" when x"8F",
		x"A1" when x"90",
		x"AF" when x"91",
		x"BD" when x"92",
		x"B3" when x"93",
		x"99" when x"94",
		x"97" when x"95",
		x"85" when x"96",
		x"8B" when x"97",
		x"D1" when x"98",
		x"DF" when x"99",
		x"CD" when x"9A",
		x"C3" when x"9B",
		x"E9" when x"9C",
		x"E7" when x"9D",
		x"F5" when x"9E",
		x"FB" when x"9F",
		x"9A" when x"A0",
		x"94" when x"A1",
		x"86" when x"A2",
		x"88" when x"A3",
		x"A2" when x"A4",
		x"AC" when x"A5",
		x"BE" when x"A6",
		x"B0" when x"A7",
		x"EA" when x"A8",
		x"E4" when x"A9",
		x"F6" when x"AA",
		x"F8" when x"AB",
		x"D2" when x"AC",
		x"DC" when x"AD",
		x"CE" when x"AE",
		x"C0" when x"AF",
		x"7A" when x"B0",
		x"74" when x"B1",
		x"66" when x"B2",
		x"68" when x"B3",
		x"42" when x"B4",
		x"4C" when x"B5",
		x"5E" when x"B6",
		x"50" when x"B7",
		x"0A" when x"B8",
		x"04" when x"B9",
		x"16" when x"BA",
		x"18" when x"BB",
		x"32" when x"BC",
		x"3C" when x"BD",
		x"2E" when x"BE",
		x"20" when x"BF",
		x"EC" when x"C0",
		x"E2" when x"C1",
		x"F0" when x"C2",
		x"FE" when x"C3",
		x"D4" when x"C4",
		x"DA" when x"C5",
		x"C8" when x"C6",
		x"C6" when x"C7",
		x"9C" when x"C8",
		x"92" when x"C9",
		x"80" when x"CA",
		x"8E" when x"CB",
		x"A4" when x"CC",
		x"AA" when x"CD",
		x"B8" when x"CE",
		x"B6" when x"CF",
		x"0C" when x"D0",
		x"02" when x"D1",
		x"10" when x"D2",
		x"1E" when x"D3",
		x"34" when x"D4",
		x"3A" when x"D5",
		x"28" when x"D6",
		x"26" when x"D7",
		x"7C" when x"D8",
		x"72" when x"D9",
		x"60" when x"DA",
		x"6E" when x"DB",
		x"44" when x"DC",
		x"4A" when x"DD",
		x"58" when x"DE",
		x"56" when x"DF",
		x"37" when x"E0",
		x"39" when x"E1",
		x"2B" when x"E2",
		x"25" when x"E3",
		x"0F" when x"E4",
		x"01" when x"E5",
		x"13" when x"E6",
		x"1D" when x"E7",
		x"47" when x"E8",
		x"49" when x"E9",
		x"5B" when x"EA",
		x"55" when x"EB",
		x"7F" when x"EC",
		x"71" when x"ED",
		x"63" when x"EE",
		x"6D" when x"EF",
		x"D7" when x"F0",
		x"D9" when x"F1",
		x"CB" when x"F2",
		x"C5" when x"F3",
		x"EF" when x"F4",
		x"E1" when x"F5",
		x"F3" when x"F6",
		x"FD" when x"F7",
		x"A7" when x"F8",
		x"A9" when x"F9",
		x"BB" when x"FA",
		x"B5" when x"FB",
		x"9F" when x"FC",
		x"91" when x"FD",
		x"83" when x"FE",
		x"8D" when x"FF",
		x"00" when others;  

end Behavioral;

